`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/05/2019 12:50:37 AM
// Design Name: 
// Module Name: bram
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module bram(
    input clk,
    input rst,
    input wena,
    input ba,
    input ha,
    input ua,
    input [7:0] addra,
    input [31:0] dina,
    output [31:0] douta
    );
    reg [7:0]mem[0:255];
    initial begin
mem[0]<=8'b00010011;
mem[1]<=8'b00000000;
mem[2]<=8'b00000000;
mem[3]<=8'b00000000;
mem[4]<=8'b10010011;
mem[5]<=8'b00000000;
mem[6]<=8'b00000000;
mem[7]<=8'b00001000;
mem[8]<=8'b00010011;
mem[9]<=8'b00000001;
mem[10]<=8'b10000000;
mem[11]<=8'b00000000;
mem[12]<=8'b10010011;
mem[13]<=8'b00000001;
mem[14]<=8'b00000000;
mem[15]<=8'b00000001;
mem[16]<=8'b00010011;
mem[17]<=8'b00000010;
mem[18]<=8'b10000000;
mem[19]<=8'b00000001;
mem[20]<=8'b10110111;
mem[21]<=8'b00010010;
mem[22]<=8'b00000000;
mem[23]<=8'b00000000;
mem[24]<=8'b00010111;
mem[25]<=8'b00010011;
mem[26]<=8'b00000000;
mem[27]<=8'b00000000;
mem[28]<=8'b00110011;
mem[29]<=8'b00000011;
mem[30]<=8'b01010011;
mem[31]<=8'b01000000;
mem[32]<=8'b10110011;
mem[33]<=8'b01110011;
mem[34]<=8'b00100010;
mem[35]<=8'b00000000;
mem[36]<=8'b01100011;
mem[37]<=8'b10001010;
mem[38]<=8'b00100011;
mem[39]<=8'b00000010;
mem[40]<=8'b10010011;
mem[41]<=8'b11010101;
mem[42]<=8'b00010101;
mem[43]<=8'b00000000;
mem[44]<=8'b01100011;
mem[45]<=8'b11010110;
mem[46]<=8'b10110110;
mem[47]<=8'b00000010;
mem[48]<=8'b01101111;
mem[49]<=8'b00000001;
mem[50]<=8'b00000000;
mem[51]<=8'b00000100;
mem[52]<=8'b00010011;
mem[53]<=8'b11010111;
mem[54]<=8'b01000110;
mem[55]<=8'b00000001;
mem[56]<=8'b10010011;
mem[57]<=8'b11010111;
mem[58]<=8'b01000101;
mem[59]<=8'b01000001;
mem[60]<=8'b00110011;
mem[61]<=8'b00101000;
mem[62]<=8'b00000111;
mem[63]<=8'b00000001;
mem[64]<=8'b01100011;
mem[65]<=8'b00000100;
mem[66]<=8'b00000101;
mem[67]<=8'b00000001;
mem[68]<=8'b01110011;
mem[69]<=8'b00000000;
mem[70]<=8'b00000000;
mem[71]<=8'b00000000;
mem[72]<=8'b00010011;
mem[73]<=8'b00000000;
mem[74]<=8'b00000000;
mem[75]<=8'b00000000;
mem[76]<=8'b00010011;
mem[77]<=8'b00000000;
mem[78]<=8'b00000000;
mem[79]<=8'b00000000;
mem[80]<=8'b00010011;
mem[81]<=8'b00000000;
mem[82]<=8'b00000000;
mem[83]<=8'b00000000;
mem[84]<=8'b01110011;
mem[85]<=8'b00000000;
mem[86]<=8'b00000000;
mem[87]<=8'b00000000;
mem[88]<=8'b00110011;
mem[89]<=8'b11100100;
mem[90]<=8'b00100001;
mem[91]<=8'b00000000;
mem[92]<=8'b10010011;
mem[93]<=8'b10010100;
mem[94]<=8'b00010001;
mem[95]<=8'b00000000;
mem[96]<=8'b00110011;
mem[97]<=8'b00110101;
mem[98]<=8'b10010100;
mem[99]<=8'b00000000;
mem[100]<=8'b10110111;
mem[101]<=8'b11110101;
mem[102]<=8'b11111111;
mem[103]<=8'b11111111;
mem[104]<=8'b10010011;
mem[105]<=8'b01100110;
mem[106]<=8'b11110000;
mem[107]<=8'b11111111;
mem[108]<=8'b11100011;
mem[109]<=8'b11111110;
mem[110]<=8'b10110110;
mem[111]<=8'b11111010;
mem[112]<=8'b00100011;
mem[113]<=8'b00000100;
mem[114]<=8'b11010000;
mem[115]<=8'b00001100;
mem[116]<=8'b10100011;
mem[117]<=8'b00010100;
mem[118]<=8'b10110000;
mem[119]<=8'b00001100;
mem[120]<=8'b10100011;
mem[121]<=8'b00100101;
mem[122]<=8'b00010000;
mem[123]<=8'b00001100;
mem[124]<=8'b10100011;
mem[125]<=8'b00010111;
mem[126]<=8'b00100000;
mem[127]<=8'b00001100;
mem[128]<=8'b00000011;
mem[129]<=8'b01000111;
mem[130]<=8'b11110000;
mem[131]<=8'b00001100;
mem[132]<=8'b01100111;
mem[133]<=8'b00000000;
mem[134]<=8'b00000111;
mem[135]<=8'b00000000;//test6

//mem[0]<=8'b00010011;
//mem[1]<=8'b00000000;
//mem[2]<=8'b00000000;
//mem[3]<=8'b00000000;  
//mem[4]<=8'b10010001;
//mem[5]<=8'b01000000;
//mem[6]<=8'b00100001;
//mem[7]<=8'b01000001;
//mem[8]<=8'b11000001;
//mem[9]<=8'b01000001;
//mem[10]<=8'b00001001;
//mem[11]<=8'b01000010;
//mem[12]<=8'b00001010;
//mem[13]<=8'b00000001;//test for compressed insts
//mem[14]<=8'b00001110;
//mem[15]<=8'b10010010;
//mem[16]<=8'b00010001;
//mem[17]<=8'b00000010;
//mem[18]<=8'b10001010;
//mem[19]<=8'b10000001;
//mem[20]<=8'b10010001;
//mem[21]<=8'b10001101;
//mem[22]<=8'b11100101;
//mem[23]<=8'b11011101;
//mem[24]<=8'b00001110;
//mem[25]<=8'b11000000;
//mem[26]<=8'b10000010;
//mem[27]<=8'b01000011;
//mem[28]<=8'b10111101;
//mem[29]<=8'b10001101;
//mem[30]<=8'b11100101;
//mem[31]<=8'b11111101;



    end
    
    always @ (posedge clk)begin
        if(wena)begin
             if(ba)begin
                mem[addra]<=dina[7:0];
            end else if(ha)begin
                mem[addra]<=dina[7:0];
                mem[addra+1]<=dina[15:8];
            end else begin
                mem[addra]<=dina[7:0];
                mem[addra+1]<=dina[15:8];
                mem[addra+2]<=dina[23:16];
                mem[addra+3]<=dina[31:24];
            end
         end
            
    end//always
  //  always @(*)begin
            assign douta={mem[addra+3],mem[addra+2], mem[addra+1], mem[addra]};
  //  end
endmodule
